////////////////////////////////////////////////////////////////////////////////
// Author: Kareem Waseem
// Course: Digital Verification using SV & UVM
//
// Description: Shift register Interface
// 
////////////////////////////////////////////////////////////////////////////////
interface sr_if ();
  logic serial_in, direction, mode;
  logic [5:0] datain, dataout;
endinterface